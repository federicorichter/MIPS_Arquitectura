module general_control #(

)
(

);

endmodule

module general_control #(
    parameter FUNC_SIZE = 6,
    parameter OP_SIZE = 6,
    parameter CONTROL_SIZE = 18
)(
    input wire [FUNC_SIZE-1:0] i_func,
    input wire [OP_SIZE-1:0] i_opcode,
    output wire [CONTROL_SIZE-1:0] o_control
);
    // TODO: Revisar los opcodes de los cases y pasar los control_reg de los comentarios a codigo xd

    // Control Bits
    localparam REG_WRITE = 0; //Reg_Write
    localparam BRANCH = 1; //Branch
    localparam UNSIGNED = 2; //Unsigned
    localparam MEM_READ = 3; //MEM_Read
    localparam MEM_WRITE = 4; //MEM_W
    localparam MASK_1 = 5; 
    localparam MASK_2 = 6;
    localparam REG_DST = 7; //Reg_dst
    localparam SHIFT_SRC = 8; //ShiftSrc
    localparam ALU_SRC = 9; //AluSrc
    localparam ALU_OP0 = 10; //Op0  (000: sub) (001: add) (010: slt) (011: and) (100: or) (101: xor) (110: lui)
    localparam ALU_OP1= 11;  //Op1
    localparam ALU_OP2 = 12; //Op2
    localparam MEM_2_REG = 13; //MEM_ToREG
    localparam J_RET_DST = 14;
    localparam EQorNE = 15;
    localparam JUMP_SRC = 16;
    localparam JUMP_OR_B = 17;

    reg [CONTROL_SIZE-1:0] control_reg;
    always @(*) begin
        casez ({i_opcode, i_func})
            // R-type instructions
            12'b000000000000: control_reg = 18'b; // SLL (shift left logical)
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 0 (shift source is rs)
            // ALU_SRC = 0 (ALU source is rt) (ALU_src)
            // ALU_OP = 111 (ALU operation is shift left logical)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b000000000010: control_reg = 18'b; // SRL
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 0 (shift source is rs)
            // ALU_SRC = 0 (ALU source is rt) (ALU_src)
            // ALU_OP = 111 (ALU operation is shift left logical)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b000000000011: control_reg = 18'b; // SRA
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 0 (shift source is rs)
            // ALU_SRC = 0 (ALU source is rt) (ALU_src)
            // ALU_OP = 111 (ALU operation is shift left logical)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b000000000100: control_reg = 18'b; // SLLV
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 1 (shift source is rs)
            // ALU_SRC = 0 (ALU source is rt) (ALU_src)
            // ALU_OP = 111 (ALU operation is shift left logical)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)            

            12'b000000000110: control_reg = 18'b; // SRLV
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 1 (shift source is rs)
            // ALU_SRC = 0 (ALU source is rt) (ALU_src)
            // ALU_OP = 111 (ALU operation is shift left logical)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)    

            12'b000000000111: control_reg = 18'b; // SRAV
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 1 (shift source is rs)
            // ALU_SRC = 0 (ALU source is rt) (ALU_src)
            // ALU_OP = 111 (ALU operation is shift left logical)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)    

            12'b000000100001: control_reg = 18'b; // ADDU
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 111 (ALU operation is add unsigned)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b000000100011: control_reg = 18'b;// SUBU
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 111 (ALU operation is add unsigned)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b000000100100: control_reg = 18'b; // AND
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 111 (ALU operation is add unsigned)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b000000100101: control_reg = 18'b; // OR
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 111 (ALU operation is add unsigned)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b000000100110: control_reg = 18'b; // XOR
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 111 (ALU operation is add unsigned)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b000000100111: control_reg = 18'b; // NOR
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 111 (ALU operation is add unsigned)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b000000101010: control_reg = 18'b; // SLT
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 111 (ALU operation is add unsigned)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b000000101011: control_reg = 18'b; // SLTU
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 1 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 111 (ALU operation is add unsigned)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            // I-type instructions
            12'b100000??????: control_reg = 18'b; // LB
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 1 (memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 1  
            // MASK_2 = 1 
            // REG_DST = 0 (destination register is rt)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is immediate)
            // ALU_OP = 001 (ALU operation is add)
            // MEM_2_REG = 1 (write memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b100001??????: control_reg = 18'b; // LH
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 1 (memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 1  
            // MASK_2 = 0  
            // REG_DST = 0 (destination register is rt)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is immediate)
            // ALU_OP = 001 (ALU operation is add)
            // MEM_2_REG = 1 (write memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)
            
            12'b100011??????: control_reg = 18'b100010010001000000; // LW
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 1 (memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0  
            // MASK_2 = 0  
            // REG_DST = 0 (destination register is rt)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is immediate)
            // ALU_OP = 001 (ALU operation is add)
            // MEM_2_REG = 1 (write memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b100111??????: control_reg = 18'b100010010001000000; // LWU
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (signed operation)
            // MEM_READ = 1 (memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0  
            // MASK_2 = 0  
            // REG_DST = 0 (destination register is rt)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is immediate)
            // ALU_OP = 001 (ALU operation is add)
            // MEM_2_REG = 1 (write memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b100100??????: control_reg = 18'b100010010001000000; // LBU
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (signed operation)
            // MEM_READ = 1 (memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 1  
            // MASK_2 = 1  
            // REG_DST = 0 (destination register is rt)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is immediate)
            // ALU_OP = 001 (ALU operation is add)
            // MEM_2_REG = 1 (write memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b100101??????: control_reg = 18'b100010010001000000; // LHU
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (signed operation)
            // MEM_READ = 1 (memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 1  
            // MASK_2 = 0  
            // REG_DST = 0 (destination register is rt)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is immediate)
            // ALU_OP = 001 (ALU operation is add)
            // MEM_2_REG = 1 (write memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b101000??????: control_reg = 18'b000000000000000000; // SB
            // REG_WRITE = 0 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (memory read)
            // MEM_WRITE = 1 (not a memory write)
            // MASK_1 = 1  
            // MASK_2 = 1  
            // REG_DST = 0 (destination register is rt)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is immediate)
            // ALU_OP = 001 (ALU operation is add)
            // MEM_2_REG = 0 (write memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b101001??????: control_reg = 18'b000000000000000000; // SH
            // REG_WRITE = 0 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (memory read)
            // MEM_WRITE = 1 (not a memory write)
            // MASK_1 = 1  
            // MASK_2 = 0  
            // REG_DST = 0 (destination register is rt)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is immediate)
            // ALU_OP = 001 (ALU operation is add)
            // MEM_2_REG = 0 (write memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b101011??????: control_reg = 18'b000000000000000000; // SW
            // REG_WRITE = 0 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (memory read)
            // MEM_WRITE = 1 (not a memory write)
            // MASK_1 = 0  
            // MASK_2 = 0  
            // REG_DST = 0 (destination register is rt)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is immediate)
            // ALU_OP = 001 (ALU operation is add)
            // MEM_2_REG = 0 (write memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b001000??????: control_reg = 18'b100001010000000000; // ADDI
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is rt)
            // ALU_OP = 001 (ALU operation is add signed)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b001001??????: control_reg = 18'b100001010000000000; // ADDIU
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is rt)
            // ALU_OP = 001 (ALU operation is add unsigned)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b001100??????: control_reg = 18'b100001010000000000; // ANDI
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is rt)
            // ALU_OP = 011 (ALU operation is and)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b001101??????: control_reg = 18'b100001010000000000; // ORI
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is rt)
            // ALU_OP = 100 (ALU operation is OR)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b001110??????: control_reg = 18'b100001010000000000; // XORI
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is rt)
            // ALU_OP = 101 (ALU operation is and)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b001111??????: control_reg = 18'b100001010000000000; // LUI
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is rt) 
            // ALU_OP = 001 (ALU operation is sum unsigned)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b001010??????: control_reg = 18'b100001010000000000; // SLTI
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is rt)
            // ALU_OP = 010 (ALU operation is slt signed)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b001011??????: control_reg = 18'b100001010000000000; // SLTIU
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 1 (unsigned operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (destination register is rd)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 1 (ALU source is rt)
            // ALU_OP = 010 (ALU operation is slt signed)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 0 (not a jump or branch instruction)

            12'b000100??????: control_reg = 18'b010000000000000000; // BEQ
            // REG_WRITE = 0 (not writing to register)
            // BRANCH = 1 (branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (not writing to register)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 000 
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 1 (branch on equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 1 (branch instruction)

            12'b000101??????: control_reg = 18'b010000000000000000; // BNE
            // REG_WRITE = 0 (not writing to register)
            // BRANCH = 1 (branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (not writing to register)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 000 
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 1 (branch on equal)
            // JUMP_SRC = 0 (not a jump instruction)
            // JUMP_OR_B = 1 (branch instruction)
            
            // J-type instructions
            12'b000010??????: control_reg = 18'b000000000000000100; // J
            // REG_WRITE = 0 (not writing to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (not writing to register)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 000 (ALU operation is add)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 0 (not a jump/return instruction)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 1 (jump instruction)
            // JUMP_OR_B = 1 (jump instruction)

            12'b000011??????: control_reg = 18'b100000000000000100; // JAL
            // Similar justificación que J, pero REG_WRITE = 1 (escribir en el registro)
            
            12'b000000??????00000: control_reg = 18'b100000000000000110; // JALR
            // REG_WRITE = 1 (write to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (not writing to register)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 000 (ALU operation is add)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 1 (es una instrucción de retorno de salto)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 1 (jump instruction)
            // JUMP_OR_B = 1 (jump instruction)

            12'b000000??????00100: control_reg = 18'b000000000000000110; // JR
            // REG_WRITE = 0 (not writing to register)
            // BRANCH = 0 (not a branch instruction)
            // UNSIGNED = 0 (signed operation)
            // MEM_READ = 0 (not a memory read)
            // MEM_WRITE = 0 (not a memory write)
            // MASK_1 = 0 (not masking)
            // MASK_2 = 0 (not masking)
            // REG_DST = 0 (not writing to register)
            // SHIFT_SRC = 0 (ALU source is rs)
            // ALU_SRC = 0 (ALU source is rt)
            // ALU_OP = 000 (ALU operation is add)
            // MEM_2_REG = 0 (not writing memory to register)
            // J_RET_DST = 1 (es una instrucción de retorno de salto)
            // EQorNE = 0 (not a branch on equal/not equal)
            // JUMP_SRC = 1 (jump instruction)
            // JUMP_OR_B = 1 (jump instruction)

            default: control_reg = 18'b000000000000000000; // Default control signals
        endcase
    end

    assign o_control = control_reg;
endmodule